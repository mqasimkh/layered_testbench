class driver;

endclass: driver